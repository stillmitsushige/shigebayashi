module template

struct Template {
	template string
}

fn parse() {}

fn execute() {}