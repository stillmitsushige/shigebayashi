/*
何も作ってない
*/

module template

struct Template {
	template string
}

fn parse(template string, target map[string]any) string {
}


fn execute() {}