module main

import commands

fn main() {
	commands.execute()
}
